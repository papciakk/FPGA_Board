use work.typedefs.all;

package model is
  constant MODEL_EDGES_NUMBER : integer := 1040;
  constant MODEL_DATA : mesh_data(1039 downto 0) := (
    X"0BCE000008360AB9FA880836",
    X"0AB9FA8808360A8BFA9C08F2",
    X"0A8BFA9C08F20B9C000008F2",
    X"0B9C000008F20BCE00000836",
    X"0A8BFA9C08F20AC1FA850931",
    X"0AC1FA8509310BD600000931",
    X"0BD6000009310B9C000008F2",
    X"0AC1FA8509310B2DFA5708F2",
    X"0B2DFA5708F20C4B000008F2",
    X"0C4B000008F20BD600000931",
    X"0B2DFA5708F20BA4FA240836",
    X"0BA4FA2408360CCD00000836",
    X"0CCD000008360C4B000008F2",
    X"0AB9FA88083607C3F61B0836",
    X"07C3F61B083607A0F63F08F2",
    X"07A0F63F08F20A8BFA9C08F2",
    X"07A0F63F08F207C9F6160931",
    X"07C9F61609310AC1FA850931",
    X"07C9F6160931081CF5C208F2",
    X"081CF5C208F20B2DFA5708F2",
    X"081CF5C208F20878F5660836",
    X"0878F56608360BA4FA240836",
    X"07C3F61B08360356F3250836",
    X"0356F32508360343F35308F2",
    X"0343F35308F207A0F63F08F2",
    X"0343F35308F20359F31E0931",
    X"0359F31E093107C9F6160931",
    X"0359F31E09310388F2B108F2",
    X"0388F2B108F2081CF5C208F2",
    X"0388F2B108F203BAF23A0836",
    X"03BAF23A08360878F5660836",
    X"0356F3250836FDDFF2110836",
    X"FDDFF2110836FDDFF24208F2",
    X"FDDFF24208F20343F35308F2",
    X"FDDFF24208F2FDDFF2090931",
    X"FDDFF20909310359F31E0931",
    X"FDDFF2090931FDDFF19308F2",
    X"FDDFF19308F20388F2B108F2",
    X"FDDFF19308F2FDDFF1120836",
    X"FDDFF112083603BAF23A0836",
    X"FDDFF2110836F806F3250836",
    X"F806F3250836F851F35308F2",
    X"F851F35308F2FDDFF24208F2",
    X"F851F35308F2F857F31E0931",
    X"F857F31E0931FDDFF2090931",
    X"F857F31E0931F834F2B108F2",
    X"F834F2B108F2FDDFF19308F2",
    X"F834F2B108F2F803F23A0836",
    X"F803F23A0836FDDFF1120836",
    X"F806F3250836F3A4F61B0836",
    X"F3A4F61B0836F3F9F63F08F2",
    X"F3F9F63F08F2F851F35308F2",
    X"F3F9F63F08F2F3E9F6160931",
    X"F3E9F6160931F857F31E0931",
    X"F3E9F6160931F39FF5C208F2",
    X"F39FF5C208F2F834F2B108F2",
    X"F39FF5C208F2F345F5660836",
    X"F345F5660836F803F23A0836",
    X"F3A4F61B0836F0E3FA880836",
    X"F0E3FA880836F124FA9C08F2",
    X"F124FA9C08F2F3F9F63F08F2",
    X"F124FA9C08F2F0F8FA850931",
    X"F0F8FA850931F3E9F6160931",
    X"F0F8FA850931F08FFA5708F2",
    X"F08FFA5708F2F39FF5C208F2",
    X"F08FFA5708F2F018FA240836",
    X"F018FA240836F345F5660836",
    X"F0E3FA880836EFEF00000836",
    X"EFEF00000836F021000008F2",
    X"F021000008F2F124FA9C08F2",
    X"F021000008F2EFE700000931",
    X"EFE700000931F0F8FA850931",
    X"EFE700000931EF72000008F2",
    X"EF72000008F2F08FFA5708F2",
    X"EF72000008F2EEF000000836",
    X"EEF000000836F018FA240836",
    X"EFEF00000836F10405780836",
    X"F10405780836F132056408F2",
    X"F132056408F2F021000008F2",
    X"F132056408F2F0FC057B0931",
    X"F0FC057B0931EFE700000931",
    X"F0FC057B0931F09005A908F2",
    X"F09005A908F2EF72000008F2",
    X"F09005A908F2F01805DC0836",
    X"F01805DC0836EEF000000836",
    X"F10405780836F3FA09E50836",
    X"F3FA09E50836F41D09C108F2",
    X"F41D09C108F2F132056408F2",
    X"F41D09C108F2F3F409EA0931",
    X"F3F409EA0931F0FC057B0931",
    X"F3F409EA0931F3A10A3E08F2",
    X"F3A10A3E08F2F09005A908F2",
    X"F3A10A3E08F2F3450A9A0836",
    X"F3450A9A0836F01805DC0836",
    X"F3FA09E50836F8670CDB0836",
    X"F8670CDB0836F87A0CAD08F2",
    X"F87A0CAD08F2F41D09C108F2",
    X"F87A0CAD08F2F8630CE20931",
    X"F8630CE20931F3F409EA0931",
    X"F8630CE20931F8350D4F08F2",
    X"F8350D4F08F2F3A10A3E08F2",
    X"F8350D4F08F2F8030DC60836",
    X"F8030DC60836F3450A9A0836",
    X"F8670CDB0836FDDF0DEF0836",
    X"FDDF0DEF0836FDDF0DBE08F2",
    X"FDDF0DBE08F2F87A0CAD08F2",
    X"FDDF0DBE08F2FDDF0DF70931",
    X"FDDF0DF70931F8630CE20931",
    X"FDDF0DF70931FDDF0E6D08F2",
    X"FDDF0E6D08F2F8350D4F08F2",
    X"FDDF0E6D08F2FDDF0EEE0836",
    X"FDDF0EEE0836F8030DC60836",
    X"FDDF0DEF083603560CDB0836",
    X"03560CDB083603430CAD08F2",
    X"03430CAD08F2FDDF0DBE08F2",
    X"03430CAD08F203590CE20931",
    X"03590CE20931FDDF0DF70931",
    X"03590CE2093103880D4F08F2",
    X"03880D4F08F2FDDF0E6D08F2",
    X"03880D4F08F203BA0DC60836",
    X"03BA0DC60836FDDF0EEE0836",
    X"03560CDB083607C309E50836",
    X"07C309E5083607A009C108F2",
    X"07A009C108F203430CAD08F2",
    X"07A009C108F207C909EA0931",
    X"07C909EA093103590CE20931",
    X"07C909EA0931081C0A3E08F2",
    X"081C0A3E08F203880D4F08F2",
    X"081C0A3E08F208780A9A0836",
    X"08780A9A083603BA0DC60836",
    X"07C309E508360AB905780836",
    X"0AB9057808360A8B056408F2",
    X"0A8B056408F207A009C108F2",
    X"0A8B056408F20AC1057B0931",
    X"0AC1057B093107C909EA0931",
    X"0AC1057B09310B2D05A908F2",
    X"0B2D05A908F2081C0A3E08F2",
    X"0B2D05A908F20BA405DC0836",
    X"0BA405DC083608780A9A0836",
    X"0AB9057808360BCE00000836",
    X"0B9C000008F20A8B056408F2",
    X"0BD6000009310AC1057B0931",
    X"0C4B000008F20B2D05A908F2",
    X"0CCD000008360BA405DC0836",
    X"0BA4FA2408360D54F96C044E",
    X"0D54F96C044E0EA10000044E",
    X"0EA10000044E0CCD00000836",
    X"0D54F96C044E0ECDF8CC0077",
    X"0ECDF8CC0077103900000077",
    X"1039000000770EA10000044E",
    X"0ECDF8CC00770FD7F85BFCC5",
    X"0FD7F85BFCC511590000FCC5",
    X"11590000FCC5103900000077",
    X"0FD7F85BFCC5103CF830F948",
    X"103CF830F94811C70000F948",
    X"11C70000F94811590000FCC5",
    X"0878F566083609C4F41A044E",
    X"09C4F41A044E0D54F96C044E",
    X"09C4F41A044E0AE6F2F80077",
    X"0AE6F2F800770ECDF8CC0077",
    X"0AE6F2F800770BB3F22BFCC5",
    X"0BB3F22BFCC50FD7F85BFCC5",
    X"0BB3F22BFCC50C01F1DEF948",
    X"0C01F1DEF948103CF830F948",
    X"03BAF23A08360472F08A044E",
    X"0472F08A044E09C4F41A044E",
    X"0472F08A044E0512EF120077",
    X"0512EF1200770AE6F2F80077",
    X"0512EF1200770584EE08FCC5",
    X"0584EE08FCC50BB3F22BFCC5",
    X"0584EE08FCC505AFEDA3F948",
    X"05AFEDA3F9480C01F1DEF948",
    X"FDDFF1120836FDDFEF3E044E",
    X"FDDFEF3E044E0472F08A044E",
    X"FDDFEF3E044EFDDFEDA60077",
    X"FDDFEDA600770512EF120077",
    X"FDDFEDA60077FDDFEC85FCC5",
    X"FDDFEC85FCC50584EE08FCC5",
    X"FDDFEC85FCC5FDDFEC18F948",
    X"FDDFEC18F94805AFEDA3F948",
    X"F803F23A0836F74BF08A044E",
    X"F74BF08A044EFDDFEF3E044E",
    X"F74BF08A044EF6ABEF120077",
    X"F6ABEF120077FDDFEDA60077",
    X"F6ABEF120077F639EE08FCC5",
    X"F639EE08FCC5FDDFEC85FCC5",
    X"F639EE08FCC5F60EEDA3F948",
    X"F60EEDA3F948FDDFEC18F948",
    X"F345F5660836F1F9F41A044E",
    X"F1F9F41A044EF74BF08A044E",
    X"F1F9F41A044EF0D7F2F80077",
    X"F0D7F2F80077F6ABEF120077",
    X"F0D7F2F80077F00AF22BFCC5",
    X"F00AF22BFCC5F639EE08FCC5",
    X"F00AF22BFCC5EFBCF1DEF948",
    X"EFBCF1DEF948F60EEDA3F948",
    X"F018FA240836EE69F96C044E",
    X"EE69F96C044EF1F9F41A044E",
    X"EE69F96C044EECF0F8CC0077",
    X"ECF0F8CC0077F0D7F2F80077",
    X"ECF0F8CC0077EBE6F85BFCC5",
    X"EBE6F85BFCC5F00AF22BFCC5",
    X"EBE6F85BFCC5EB81F830F948",
    X"EB81F830F948EFBCF1DEF948",
    X"EEF000000836ED1C0000044E",
    X"ED1C0000044EEE69F96C044E",
    X"ED1C0000044EEB8400000077",
    X"EB8400000077ECF0F8CC0077",
    X"EB8400000077EA630000FCC5",
    X"EA630000FCC5EBE6F85BFCC5",
    X"EA630000FCC5E9F60000F948",
    X"E9F60000F948EB81F830F948",
    X"F01805DC0836EE690694044E",
    X"EE690694044EED1C0000044E",
    X"EE690694044EECF007340077",
    X"ECF007340077EB8400000077",
    X"ECF007340077EBE607A5FCC5",
    X"EBE607A5FCC5EA630000FCC5",
    X"EBE607A5FCC5EB8107D0F948",
    X"EB8107D0F948E9F60000F948",
    X"F3450A9A0836F1F90BE6044E",
    X"F1F90BE6044EEE690694044E",
    X"F1F90BE6044EF0D70D080077",
    X"F0D70D080077ECF007340077",
    X"F0D70D080077F00A0DD5FCC5",
    X"F00A0DD5FCC5EBE607A5FCC5",
    X"F00A0DD5FCC5EFBC0E22F948",
    X"EFBC0E22F948EB8107D0F948",
    X"F8030DC60836F74B0F76044E",
    X"F74B0F76044EF1F90BE6044E",
    X"F74B0F76044EF6AB10EE0077",
    X"F6AB10EE0077F0D70D080077",
    X"F6AB10EE0077F63911F8FCC5",
    X"F63911F8FCC5F00A0DD5FCC5",
    X"F63911F8FCC5F60E125DF948",
    X"F60E125DF948EFBC0E22F948",
    X"FDDF0EEE0836FDDF10C2044E",
    X"FDDF10C2044EF74B0F76044E",
    X"FDDF10C2044EFDDF125A0077",
    X"FDDF125A0077F6AB10EE0077",
    X"FDDF125A0077FDDF137BFCC5",
    X"FDDF137BFCC5F63911F8FCC5",
    X"FDDF137BFCC5FDDF13E8F948",
    X"FDDF13E8F948F60E125DF948",
    X"03BA0DC6083604720F76044E",
    X"04720F76044EFDDF10C2044E",
    X"04720F76044E051210EE0077",
    X"051210EE0077FDDF125A0077",
    X"051210EE0077058411F8FCC5",
    X"058411F8FCC5FDDF137BFCC5",
    X"058411F8FCC505AF125DF948",
    X"05AF125DF948FDDF13E8F948",
    X"08780A9A083609C40BE6044E",
    X"09C40BE6044E04720F76044E",
    X"09C40BE6044E0AE60D080077",
    X"0AE60D080077051210EE0077",
    X"0AE60D0800770BB30DD5FCC5",
    X"0BB30DD5FCC5058411F8FCC5",
    X"0BB30DD5FCC50C010E22F948",
    X"0C010E22F94805AF125DF948",
    X"0BA405DC08360D540694044E",
    X"0D540694044E09C40BE6044E",
    X"0D540694044E0ECD07340077",
    X"0ECD073400770AE60D080077",
    X"0ECD073400770FD707A5FCC5",
    X"0FD707A5FCC50BB30DD5FCC5",
    X"0FD707A5FCC5103C07D0F948",
    X"103C07D0F9480C010E22F948",
    X"0EA10000044E0D540694044E",
    X"1039000000770ECD07340077",
    X"11590000FCC50FD707A5FCC5",
    X"11C70000F948103C07D0F948",
    X"103CF830F9480F84F87EF655",
    X"0F84F87EF65511000000F655",
    X"11000000F65511C70000F948",
    X"0F84F87EF6550DF0F92AF426",
    X"0DF0F92AF4260F4A0000F426",
    X"0F4A0000F42611000000F655",
    X"0DF0F92AF4260C5CF9D6F2AB",
    X"0C5CF9D6F2AB0D940000F2AB",
    X"0D940000F2AB0F4A0000F426",
    X"0C5CF9D6F2AB0BA4FA24F1D1",
    X"0BA4FA24F1D10CCD0000F1D1",
    X"0CCD0000F1D10D940000F2AB",
    X"0C01F1DEF9480B73F26BF655",
    X"0B73F26BF6550F84F87EF655",
    X"0B73F26BF6550A3CF3A2F426",
    X"0A3CF3A2F4260DF0F92AF426",
    X"0A3CF3A2F4260905F4D9F2AB",
    X"0905F4D9F2AB0C5CF9D6F2AB",
    X"0905F4D9F2AB0878F566F1D1",
    X"0878F566F1D10BA4FA24F1D1",
    X"05AFEDA3F9480560EE5AF655",
    X"0560EE5AF6550B73F26BF655",
    X"0560EE5AF65504B4EFEEF426",
    X"04B4EFEEF4260A3CF3A2F426",
    X"04B4EFEEF4260409F182F2AB",
    X"0409F182F2AB0905F4D9F2AB",
    X"0409F182F2AB03BAF23AF1D1",
    X"03BAF23AF1D10878F566F1D1",
    X"FDDFEC18F948FDDFECDFF655",
    X"FDDFECDFF6550560EE5AF655",
    X"FDDFECDFF655FDDFEE95F426",
    X"FDDFEE95F42604B4EFEEF426",
    X"FDDFEE95F426FDDFF04BF2AB",
    X"FDDFF04BF2AB0409F182F2AB",
    X"FDDFF04BF2ABFDDFF112F1D1",
    X"FDDFF112F1D103BAF23AF1D1",
    X"F60EEDA3F948F65DEE5AF655",
    X"F65DEE5AF655FDDFECDFF655",
    X"F65DEE5AF655F708EFEEF426",
    X"F708EFEEF426FDDFEE95F426",
    X"F708EFEEF426F7B4F182F2AB",
    X"F7B4F182F2ABFDDFF04BF2AB",
    X"F7B4F182F2ABF803F23AF1D1",
    X"F803F23AF1D1FDDFF112F1D1",
    X"EFBCF1DEF948F049F26BF655",
    X"F049F26BF655F65DEE5AF655",
    X"F049F26BF655F180F3A2F426",
    X"F180F3A2F426F708EFEEF426",
    X"F180F3A2F426F2B7F4D9F2AB",
    X"F2B7F4D9F2ABF7B4F182F2AB",
    X"F2B7F4D9F2ABF345F566F1D1",
    X"F345F566F1D1F803F23AF1D1",
    X"EB81F830F948EC39F87EF655",
    X"EC39F87EF655F049F26BF655",
    X"EC39F87EF655EDCDF92AF426",
    X"EDCDF92AF426F180F3A2F426",
    X"EDCDF92AF426EF61F9D6F2AB",
    X"EF61F9D6F2ABF2B7F4D9F2AB",
    X"EF61F9D6F2ABF018FA24F1D1",
    X"F018FA24F1D1F345F566F1D1",
    X"E9F60000F948EABD0000F655",
    X"EABD0000F655EC39F87EF655",
    X"EABD0000F655EC730000F426",
    X"EC730000F426EDCDF92AF426",
    X"EC730000F426EE290000F2AB",
    X"EE290000F2ABEF61F9D6F2AB",
    X"EE290000F2ABEEF00000F1D1",
    X"EEF00000F1D1F018FA24F1D1",
    X"EB8107D0F948EC390782F655",
    X"EC390782F655EABD0000F655",
    X"EC390782F655EDCD06D6F426",
    X"EDCD06D6F426EC730000F426",
    X"EDCD06D6F426EF61062AF2AB",
    X"EF61062AF2ABEE290000F2AB",
    X"EF61062AF2ABF01805DCF1D1",
    X"F01805DCF1D1EEF00000F1D1",
    X"EFBC0E22F948F0490D95F655",
    X"F0490D95F655EC390782F655",
    X"F0490D95F655F1800C5EF426",
    X"F1800C5EF426EDCD06D6F426",
    X"F1800C5EF426F2B70B27F2AB",
    X"F2B70B27F2ABEF61062AF2AB",
    X"F2B70B27F2ABF3450A9AF1D1",
    X"F3450A9AF1D1F01805DCF1D1",
    X"F60E125DF948F65D11A6F655",
    X"F65D11A6F655F0490D95F655",
    X"F65D11A6F655F7081012F426",
    X"F7081012F426F1800C5EF426",
    X"F7081012F426F7B40E7EF2AB",
    X"F7B40E7EF2ABF2B70B27F2AB",
    X"F7B40E7EF2ABF8030DC6F1D1",
    X"F8030DC6F1D1F3450A9AF1D1",
    X"FDDF13E8F948FDDF1321F655",
    X"FDDF1321F655F65D11A6F655",
    X"FDDF1321F655FDDF116BF426",
    X"FDDF116BF426F7081012F426",
    X"FDDF116BF426FDDF0FB5F2AB",
    X"FDDF0FB5F2ABF7B40E7EF2AB",
    X"FDDF0FB5F2ABFDDF0EEEF1D1",
    X"FDDF0EEEF1D1F8030DC6F1D1",
    X"05AF125DF948056011A6F655",
    X"056011A6F655FDDF1321F655",
    X"056011A6F65504B41012F426",
    X"04B41012F426FDDF116BF426",
    X"04B41012F42604090E7EF2AB",
    X"04090E7EF2ABFDDF0FB5F2AB",
    X"04090E7EF2AB03BA0DC6F1D1",
    X"03BA0DC6F1D1FDDF0EEEF1D1",
    X"0C010E22F9480B730D95F655",
    X"0B730D95F655056011A6F655",
    X"0B730D95F6550A3C0C5EF426",
    X"0A3C0C5EF42604B41012F426",
    X"0A3C0C5EF42609050B27F2AB",
    X"09050B27F2AB04090E7EF2AB",
    X"09050B27F2AB08780A9AF1D1",
    X"08780A9AF1D103BA0DC6F1D1",
    X"103C07D0F9480F840782F655",
    X"0F840782F6550B730D95F655",
    X"0F840782F6550DF006D6F426",
    X"0DF006D6F4260A3C0C5EF426",
    X"0DF006D6F4260C5C062AF2AB",
    X"0C5C062AF2AB09050B27F2AB",
    X"0C5C062AF2AB0BA405DCF1D1",
    X"0BA405DCF1D108780A9AF1D1",
    X"11000000F6550F840782F655",
    X"0F4A0000F4260DF006D6F426",
    X"0D940000F2AB0C5C062AF2AB",
    X"0CCD0000F1D10BA405DCF1D1",
    X"0BA4FA24F1D10B55FA46F145",
    X"0B55FA46F1450C760000F145",
    X"0C760000F1450CCD0000F1D1",
    X"0B55FA46F14509AAFAFCF0CA",
    X"09AAFAFCF0CA0AA70000F0CA",
    X"0AA70000F0CA0C760000F145",
    X"09AAFAFCF0CA058AFCBDF073",
    X"058AFCBDF073062F0000F073",
    X"062F0000F0730AA70000F0CA",
    X"058AFCBDF073FDDF0000F053",
    X"FDDF0000F053062F0000F073",
    X"0878F566F1D1083BF5A4F145",
    X"083BF5A4F1450B55FA46F145",
    X"083BF5A4F14506F2F6EDF0CA",
    X"06F2F6EDF0CA09AAFAFCF0CA",
    X"06F2F6EDF0CA03C6FA19F073",
    X"03C6FA19F073058AFCBDF073",
    X"03C6FA19F073FDDF0000F053",
    X"03BAF23AF1D10398F28AF145",
    X"0398F28AF145083BF5A4F145",
    X"0398F28AF14502E3F435F0CA",
    X"02E3F435F0CA06F2F6EDF0CA",
    X"02E3F435F0CA0122F854F073",
    X"0122F854F07303C6FA19F073",
    X"0122F854F073FDDF0000F053",
    X"FDDFF112F1D1FDDFF168F145",
    X"FDDFF168F1450398F28AF145",
    X"FDDFF168F145FDDFF337F0CA",
    X"FDDFF337F0CA02E3F435F0CA",
    X"FDDFF337F0CAFDDFF7AFF073",
    X"FDDFF7AFF0730122F854F073",
    X"FDDFF7AFF073FDDF0000F053",
    X"F803F23AF1D1F825F28AF145",
    X"F825F28AF145FDDFF168F145",
    X"F825F28AF145F8DAF435F0CA",
    X"F8DAF435F0CAFDDFF337F0CA",
    X"F8DAF435F0CAFA9BF854F073",
    X"FA9BF854F073FDDFF7AFF073",
    X"FA9BF854F073FDDF0000F053",
    X"F345F566F1D1F382F5A4F145",
    X"F382F5A4F145F825F28AF145",
    X"F382F5A4F145F4CBF6EDF0CA",
    X"F4CBF6EDF0CAF8DAF435F0CA",
    X"F4CBF6EDF0CAF7F7FA19F073",
    X"F7F7FA19F073FA9BF854F073",
    X"F7F7FA19F073FDDF0000F053",
    X"F018FA24F1D1F068FA46F145",
    X"F068FA46F145F382F5A4F145",
    X"F068FA46F145F213FAFCF0CA",
    X"F213FAFCF0CAF4CBF6EDF0CA",
    X"F213FAFCF0CAF633FCBDF073",
    X"F633FCBDF073F7F7FA19F073",
    X"F633FCBDF073FDDF0000F053",
    X"EEF00000F1D1EF470000F145",
    X"EF470000F145F068FA46F145",
    X"EF470000F145F1160000F0CA",
    X"F1160000F0CAF213FAFCF0CA",
    X"F1160000F0CAF58E0000F073",
    X"F58E0000F073F633FCBDF073",
    X"F58E0000F073FDDF0000F053",
    X"F01805DCF1D1F06805BAF145",
    X"F06805BAF145EF470000F145",
    X"F06805BAF145F2130504F0CA",
    X"F2130504F0CAF1160000F0CA",
    X"F2130504F0CAF6330343F073",
    X"F6330343F073F58E0000F073",
    X"F6330343F073FDDF0000F053",
    X"F3450A9AF1D1F3820A5CF145",
    X"F3820A5CF145F06805BAF145",
    X"F3820A5CF145F4CB0913F0CA",
    X"F4CB0913F0CAF2130504F0CA",
    X"F4CB0913F0CAF7F705E7F073",
    X"F7F705E7F073F6330343F073",
    X"F7F705E7F073FDDF0000F053",
    X"F8030DC6F1D1F8250D76F145",
    X"F8250D76F145F3820A5CF145",
    X"F8250D76F145F8DA0BCBF0CA",
    X"F8DA0BCBF0CAF4CB0913F0CA",
    X"F8DA0BCBF0CAFA9B07ACF073",
    X"FA9B07ACF073F7F705E7F073",
    X"FA9B07ACF073FDDF0000F053",
    X"FDDF0EEEF1D1FDDF0E98F145",
    X"FDDF0E98F145F8250D76F145",
    X"FDDF0E98F145FDDF0CC9F0CA",
    X"FDDF0CC9F0CAF8DA0BCBF0CA",
    X"FDDF0CC9F0CAFDDF0851F073",
    X"FDDF0851F073FA9B07ACF073",
    X"FDDF0851F073FDDF0000F053",
    X"03BA0DC6F1D103980D76F145",
    X"03980D76F145FDDF0E98F145",
    X"03980D76F14502E30BCBF0CA",
    X"02E30BCBF0CAFDDF0CC9F0CA",
    X"02E30BCBF0CA012207ACF073",
    X"012207ACF073FDDF0851F073",
    X"012207ACF073FDDF0000F053",
    X"08780A9AF1D1083B0A5CF145",
    X"083B0A5CF14503980D76F145",
    X"083B0A5CF14506F20913F0CA",
    X"06F20913F0CA02E30BCBF0CA",
    X"06F20913F0CA03C605E7F073",
    X"03C605E7F073012207ACF073",
    X"03C605E7F073FDDF0000F053",
    X"0BA405DCF1D10B5505BAF145",
    X"0B5505BAF145083B0A5CF145",
    X"0B5505BAF14509AA0504F0CA",
    X"09AA0504F0CA06F20913F0CA",
    X"09AA0504F0CA058A0343F073",
    X"058A0343F07303C605E7F073",
    X"058A0343F073FDDF0000F053",
    X"0C760000F1450B5505BAF145",
    X"0AA70000F0CA09AA0504F0CA",
    X"062F0000F073058A0343F073",
    X"EDF10000047AEE19FE5204D4",
    X"EE19FE5204D4E927FE5204CA",
    X"E927FE5204CAE94B00000471",
    X"E94B00000471EDF10000047A",
    X"E927FE5204CAE586FE520481",
    X"E586FE520481E5DB00000433",
    X"E5DB00000433E94B00000471",
    X"E586FE520481E34AFE5203BC",
    X"E34AFE5203BCE3B900000388",
    X"E3B900000388E5DB00000433",
    X"E34AFE5203BCE287FE52023D",
    X"E287FE52023DE2FE0000023D",
    X"E2FE0000023DE3B900000388",
    X"EE19FE5204D4EE71FDC30599",
    X"EE71FDC30599E8D9FDC3058C",
    X"E8D9FDC3058CE927FE5204CA",
    X"E8D9FDC3058CE4CCFDC3052E",
    X"E4CCFDC3052EE586FE520481",
    X"E4CCFDC3052EE255FDC3042E",
    X"E255FDC3042EE34AFE5203BC",
    X"E255FDC3042EE180FDC3023D",
    X"E180FDC3023DE287FE52023D",
    X"EE71FDC30599EEC8FE52065E",
    X"EEC8FE52065EE88BFE52064E",
    X"E88BFE52064EE8D9FDC3058C",
    X"E88BFE52064EE412FE5205DA",
    X"E412FE5205DAE4CCFDC3052E",
    X"E412FE5205DAE160FE5204A0",
    X"E160FE5204A0E255FDC3042E",
    X"E160FE5204A0E079FE52023D",
    X"E079FE52023DE180FDC3023D",
    X"EEC8FE52065EEEF0000006B8",
    X"EEF0000006B8E868000006A6",
    X"E868000006A6E88BFE52064E",
    X"E868000006A6E3BD00000628",
    X"E3BD00000628E412FE5205DA",
    X"E3BD00000628E0F0000004D4",
    X"E0F0000004D4E160FE5204A0",
    X"E0F0000004D4E0020000023D",
    X"E0020000023DE079FE52023D",
    X"EEF0000006B8EEC801AE065E",
    X"EEC801AE065EE88B01AE064E",
    X"E88B01AE064EE868000006A6",
    X"E88B01AE064EE41201AE05DA",
    X"E41201AE05DAE3BD00000628",
    X"E41201AE05DAE16001AE04A0",
    X"E16001AE04A0E0F0000004D4",
    X"E16001AE04A0E07901AE023D",
    X"E07901AE023DE0020000023D",
    X"EEC801AE065EEE71023D0599",
    X"EE71023D0599E8D9023D058C",
    X"E8D9023D058CE88B01AE064E",
    X"E8D9023D058CE4CC023D052E",
    X"E4CC023D052EE41201AE05DA",
    X"E4CC023D052EE255023D042E",
    X"E255023D042EE16001AE04A0",
    X"E255023D042EE180023D023D",
    X"E180023D023DE07901AE023D",
    X"EE71023D0599EE1901AE04D4",
    X"EE1901AE04D4E92701AE04CA",
    X"E92701AE04CAE8D9023D058C",
    X"E92701AE04CAE58601AE0481",
    X"E58601AE0481E4CC023D052E",
    X"E58601AE0481E34A01AE03BC",
    X"E34A01AE03BCE255023D042E",
    X"E34A01AE03BCE28701AE023D",
    X"E28701AE023DE180023D023D",
    X"EE1901AE04D4EDF10000047A",
    X"E94B00000471E92701AE04CA",
    X"E5DB00000433E58601AE0481",
    X"E3B900000388E34A01AE03BC",
    X"E2FE0000023DE28701AE023D",
    X"E287FE52023DE2F5FE520003",
    X"E2F5FE520003E36200000035",
    X"E36200000035E2FE0000023D",
    X"E2F5FE520003E44FFE52FD77",
    X"E44FFE52FD77E49C0000FDC3",
    X"E49C0000FDC3E36200000035",
    X"E44FFE52FD77E6ABFE52FAF1",
    X"E6ABFE52FAF1E6C60000FB50",
    X"E6C60000FB50E49C0000FDC3",
    X"E6ABFE52FAF1EA1EFE52F8D1",
    X"EA1EFE52F8D1E9F60000F948",
    X"E9F60000F948E6C60000FB50",
    X"E180FDC3023DE206FDC3FF96",
    X"E206FDC3FF96E2F5FE520003",
    X"E206FDC3FF96E3A5FDC3FCCE",
    X"E3A5FDC3FCCEE44FFE52FD77",
    X"E3A5FDC3FCCEE66FFDC3FA22",
    X"E66FFDC3FA22E6ABFE52FAF1",
    X"E66FFDC3FA22EA75FDC3F7CA",
    X"EA75FDC3F7CAEA1EFE52F8D1",
    X"E079FE52023DE117FE52FF27",
    X"E117FE52FF27E206FDC3FF96",
    X"E117FE52FF27E2FCFE52FC26",
    X"E2FCFE52FC26E3A5FDC3FCCE",
    X"E2FCFE52FC26E634FE52F952",
    X"E634FE52F952E66FFDC3FA22",
    X"E634FE52F952EACDFE52F6C3",
    X"EACDFE52F6C3EA75FDC3F7CA",
    X"E0020000023DE0AB0000FEF5",
    X"E0AB0000FEF5E117FE52FF27",
    X"E0AB0000FEF5E2AE0000FBD9",
    X"E2AE0000FBD9E2FCFE52FC26",
    X"E2AE0000FBD9E6180000F8F3",
    X"E6180000F8F3E634FE52F952",
    X"E6180000F8F3EAF50000F64C",
    X"EAF50000F64CEACDFE52F6C3",
    X"E07901AE023DE11701AEFF27",
    X"E11701AEFF27E0AB0000FEF5",
    X"E11701AEFF27E2FC01AEFC26",
    X"E2FC01AEFC26E2AE0000FBD9",
    X"E2FC01AEFC26E63401AEF952",
    X"E63401AEF952E6180000F8F3",
    X"E63401AEF952EACD01AEF6C3",
    X"EACD01AEF6C3EAF50000F64C",
    X"E180023D023DE206023DFF96",
    X"E206023DFF96E11701AEFF27",
    X"E206023DFF96E3A5023DFCCE",
    X"E3A5023DFCCEE2FC01AEFC26",
    X"E3A5023DFCCEE66F023DFA22",
    X"E66F023DFA22E63401AEF952",
    X"E66F023DFA22EA75023DF7CA",
    X"EA75023DF7CAEACD01AEF6C3",
    X"E28701AE023DE2F501AE0003",
    X"E2F501AE0003E206023DFF96",
    X"E2F501AE0003E44F01AEFD77",
    X"E44F01AEFD77E3A5023DFCCE",
    X"E44F01AEFD77E6AB01AEFAF1",
    X"E6AB01AEFAF1E66F023DFA22",
    X"E6AB01AEFAF1EA1E01AEF8D1",
    X"EA1E01AEF8D1EA75023DF7CA",
    X"E36200000035E2F501AE0003",
    X"E49C0000FDC3E44F01AEFD77",
    X"E6C60000FB50E6AB01AEFAF1",
    X"E9F60000F948EA1E01AEF8D1",
    X"0ECA0000FE820ECAFC4EFD3A",
    X"0ECAFC4EFD3A13EEFCAAFEA7",
    X"13EEFCAAFEA713910000FF9B",
    X"13910000FF9B0ECA0000FE82",
    X"13EEFCAAFEA7161AFD7401AF",
    X"161AFD7401AF15A20000023D",
    X"15A20000023D13910000FF9B",
    X"161AFD7401AF1757FE3E053C",
    X"1757FE3E053C16C50000056F",
    X"16C50000056F15A20000023D",
    X"1757FE3E053C19AEFE9A0836",
    X"19AEFE9A083618BF00000836",
    X"18BF0000083616C50000056F",
    X"0ECAFC4EFD3A0ECAFB13FA67",
    X"0ECAFB13FA6714BCFB8DFC8F",
    X"14BCFB8DFC8F13EEFCAAFEA7",
    X"14BCFB8DFC8F1721FC9B0077",
    X"1721FC9B0077161AFD7401AF",
    X"1721FC9B00771897FDA804CB",
    X"1897FDA804CB1757FE3E053C",
    X"1897FDA804CB1BBBFE230836",
    X"1BBBFE23083619AEFE9A0836",
    X"0ECAFB13FA670ECAFC4EF794",
    X"0ECAFC4EF7941589FCAAFA78",
    X"1589FCAAFA7814BCFB8DFC8F",
    X"1589FCAAFA781828FD74FF40",
    X"1828FD74FF401721FC9B0077",
    X"1828FD74FF4019D7FE3E045A",
    X"19D7FE3E045A1897FDA804CB",
    X"19D7FE3E045A1DC9FE9A0836",
    X"1DC9FE9A08361BBBFE230836",
    X"0ECAFC4EF7940ECA0000F64C",
    X"0ECA0000F64C15E60000F984",
    X"15E60000F9841589FCAAFA78",
    X"15E60000F984189F0000FEB2",
    X"189F0000FEB21828FD74FF40",
    X"189F0000FEB21A6900000427",
    X"1A690000042719D7FE3E045A",
    X"1A69000004271EB800000836",
    X"1EB8000008361DC9FE9A0836",
    X"0ECA0000F64C0ECA03B2F794",
    X"0ECA03B2F79415890356FA78",
    X"15890356FA7815E60000F984",
    X"15890356FA781828028CFF40",
    X"1828028CFF40189F0000FEB2",
    X"1828028CFF4019D701C2045A",
    X"19D701C2045A1A6900000427",
    X"19D701C2045A1DC901660836",
    X"1DC9016608361EB800000836",
    X"0ECA03B2F7940ECA04EDFA67",
    X"0ECA04EDFA6714BC0473FC8F",
    X"14BC0473FC8F15890356FA78",
    X"14BC0473FC8F172103650077",
    X"1721036500771828028CFF40",
    X"1721036500771897025804CB",
    X"1897025804CB19D701C2045A",
    X"1897025804CB1BBB01DD0836",
    X"1BBB01DD08361DC901660836",
    X"0ECA04EDFA670ECA03B2FD3A",
    X"0ECA03B2FD3A13EE0356FEA7",
    X"13EE0356FEA714BC0473FC8F",
    X"13EE0356FEA7161A028C01AF",
    X"161A028C01AF172103650077",
    X"161A028C01AF175701C2053C",
    X"175701C2053C1897025804CB",
    X"175701C2053C19AE01660836",
    X"19AE016608361BBB01DD0836",
    X"0ECA03B2FD3A0ECA0000FE82",
    X"13910000FF9B13EE0356FEA7",
    X"15A20000023D161A028C01AF",
    X"16C50000056F175701C2053C",
    X"18BF0000083619AE01660836",
    X"19AEFE9A08361A76FEB108A7",
    X"1A76FEB108A71976000008A2",
    X"1976000008A218BF00000836",
    X"1A76FEB108A71AEEFEE208CE",
    X"1AEEFEE208CE19FD000008C5",
    X"19FD000008C51976000008A2",
    X"1AEEFEE208CE1AF1FF1308A9",
    X"1AF1FF1308A91A25000008A2",
    X"1A25000008A219FD000008C5",
    X"1AF1FF1308A91A5DFF290836",
    X"1A5DFF29083619BE00000836",
    X"19BE000008361A25000008A2",
    X"1BBBFE2308361CA9FE4108B2",
    X"1CA9FE4108B21A76FEB108A7",
    X"1CA9FE4108B21CFEFE8208E0",
    X"1CFEFE8208E01AEEFEE208CE",
    X"1CFEFE8208E01CB2FEC408B9",
    X"1CB2FEC408B91AF1FF1308A9",
    X"1CB2FEC408B91BBBFEE20836",
    X"1BBBFEE208361A5DFF290836",
    X"1DC9FE9A08361EDCFEB108BE",
    X"1EDCFEB108BE1CA9FE4108B2",
    X"1EDCFEB108BE1F0EFEE208F3",
    X"1F0EFEE208F31CFEFE8208E0",
    X"1F0EFEE208F31E72FF1308C9",
    X"1E72FF1308C91CB2FEC408B9",
    X"1E72FF1308C91D1AFF290836",
    X"1D1AFF2908361BBBFEE20836",
    X"1EB8000008361FDC000008C3",
    X"1FDC000008C31EDCFEB108BE",
    X"1FDC000008C31FFE000008FB",
    X"1FFE000008FB1F0EFEE208F3",
    X"1FFE000008FB1F3E000008D1",
    X"1F3E000008D11E72FF1308C9",
    X"1F3E000008D11DB900000836",
    X"1DB9000008361D1AFF290836",
    X"1DC9016608361EDC014F08BE",
    X"1EDC014F08BE1FDC000008C3",
    X"1EDC014F08BE1F0E011E08F3",
    X"1F0E011E08F31FFE000008FB",
    X"1F0E011E08F31E7200ED08C9",
    X"1E7200ED08C91F3E000008D1",
    X"1E7200ED08C91D1A00D70836",
    X"1D1A00D708361DB900000836",
    X"1BBB01DD08361CA901BF08B2",
    X"1CA901BF08B21EDC014F08BE",
    X"1CA901BF08B21CFE017E08E0",
    X"1CFE017E08E01F0E011E08F3",
    X"1CFE017E08E01CB2013C08B9",
    X"1CB2013C08B91E7200ED08C9",
    X"1CB2013C08B91BBB011E0836",
    X"1BBB011E08361D1A00D70836",
    X"19AE016608361A76014F08A7",
    X"1A76014F08A71CA901BF08B2",
    X"1A76014F08A71AEE011E08CE",
    X"1AEE011E08CE1CFE017E08E0",
    X"1AEE011E08CE1AF100ED08A9",
    X"1AF100ED08A91CB2013C08B9",
    X"1AF100ED08A91A5D00D70836",
    X"1A5D00D708361BBB011E0836",
    X"1976000008A21A76014F08A7",
    X"19FD000008C51AEE011E08CE",
    X"1A25000008A21AF100ED08A9",
    X"19BE000008361A5D00D70836",
    X"00FFFEAB0F30014200000F30",
    X"014200000F30FDDF00000FAD",
    X"FDDF00000FAD00FFFEAB0F30",
    X"00FFFEAB0F3000DAFEBB0DFF",
    X"00DAFEBB0DFF011A00000DFF",
    X"011A00000DFF014200000F30",
    X"00DAFEBB0DFFFFAEFF3B0C87",
    X"FFAEFF3B0C87FFD500000C87",
    X"FFD500000C87011A00000DFF",
    X"FFAEFF3B0C87FFB5FF380B33",
    X"FFB5FF380B33FFDD00000B33",
    X"FFDD00000B33FFD500000C87",
    X"0047FD970F3000FFFEAB0F30",
    X"FDDF00000FAD0047FD970F30",
    X"0047FD970F30002BFDB40DFF",
    X"002BFDB40DFF00DAFEBB0DFF",
    X"002BFDB40DFFFF43FE9C0C87",
    X"FF43FE9C0C87FFAEFF3B0C87",
    X"FF43FE9C0C87FF49FE970B33",
    X"FF49FE970B33FFB5FF380B33",
    X"FF35FCDF0F300047FD970F30",
    X"FDDF00000FADFF35FCDF0F30",
    X"FF35FCDF0F30FF25FD040DFF",
    X"FF25FD040DFF002BFDB40DFF",
    X"FF25FD040DFFFEA4FE320C87",
    X"FEA4FE320C87FF43FE9C0C87",
    X"FEA4FE320C87FEA7FE2A0B33",
    X"FEA7FE2A0B33FF49FE970B33",
    X"FDDFFC9C0F30FF35FCDF0F30",
    X"FDDF00000FADFDDFFC9C0F30",
    X"FDDFFC9C0F30FDDFFCC40DFF",
    X"FDDFFCC40DFFFF25FD040DFF",
    X"FDDFFCC40DFFFDDFFE0B0C87",
    X"FDDFFE0B0C87FEA4FE320C87",
    X"FDDFFE0B0C87FDDFFE030B33",
    X"FDDFFE030B33FEA7FE2A0B33",
    X"FC89FCDF0F30FDDFFC9C0F30",
    X"FDDF00000FADFC89FCDF0F30",
    X"FC89FCDF0F30FC99FD040DFF",
    X"FC99FD040DFFFDDFFCC40DFF",
    X"FC99FD040DFFFD1AFE320C87",
    X"FD1AFE320C87FDDFFE0B0C87",
    X"FD1AFE320C87FD17FE2A0B33",
    X"FD17FE2A0B33FDDFFE030B33",
    X"FB76FD970F30FC89FCDF0F30",
    X"FDDF00000FADFB76FD970F30",
    X"FB76FD970F30FB92FDB40DFF",
    X"FB92FDB40DFFFC99FD040DFF",
    X"FB92FDB40DFFFC7AFE9C0C87",
    X"FC7AFE9C0C87FD1AFE320C87",
    X"FC7AFE9C0C87FC75FE970B33",
    X"FC75FE970B33FD17FE2A0B33",
    X"FABEFEAB0F30FB76FD970F30",
    X"FDDF00000FADFABEFEAB0F30",
    X"FABEFEAB0F30FAE3FEBB0DFF",
    X"FAE3FEBB0DFFFB92FDB40DFF",
    X"FAE3FEBB0DFFFC10FF3B0C87",
    X"FC10FF3B0C87FC7AFE9C0C87",
    X"FC10FF3B0C87FC09FF380B33",
    X"FC09FF380B33FC75FE970B33",
    X"FA7B00000F30FABEFEAB0F30",
    X"FDDF00000FADFA7B00000F30",
    X"FA7B00000F30FAA300000DFF",
    X"FAA300000DFFFAE3FEBB0DFF",
    X"FAA300000DFFFBE900000C87",
    X"FBE900000C87FC10FF3B0C87",
    X"FBE900000C87FBE100000B33",
    X"FBE100000B33FC09FF380B33",
    X"FABE01550F30FA7B00000F30",
    X"FDDF00000FADFABE01550F30",
    X"FABE01550F30FAE301450DFF",
    X"FAE301450DFFFAA300000DFF",
    X"FAE301450DFFFC1000C50C87",
    X"FC1000C50C87FBE900000C87",
    X"FC1000C50C87FC0900C80B33",
    X"FC0900C80B33FBE100000B33",
    X"FB7602690F30FABE01550F30",
    X"FDDF00000FADFB7602690F30",
    X"FB7602690F30FB92024C0DFF",
    X"FB92024C0DFFFAE301450DFF",
    X"FB92024C0DFFFC7A01640C87",
    X"FC7A01640C87FC1000C50C87",
    X"FC7A01640C87FC7501690B33",
    X"FC7501690B33FC0900C80B33",
    X"FC8903210F30FB7602690F30",
    X"FDDF00000FADFC8903210F30",
    X"FC8903210F30FC9902FC0DFF",
    X"FC9902FC0DFFFB92024C0DFF",
    X"FC9902FC0DFFFD1A01CE0C87",
    X"FD1A01CE0C87FC7A01640C87",
    X"FD1A01CE0C87FD1701D60B33",
    X"FD1701D60B33FC7501690B33",
    X"FDDF03640F30FC8903210F30",
    X"FDDF00000FADFDDF03640F30",
    X"FDDF03640F30FDDF033C0DFF",
    X"FDDF033C0DFFFC9902FC0DFF",
    X"FDDF033C0DFFFDDF01F50C87",
    X"FDDF01F50C87FD1A01CE0C87",
    X"FDDF01F50C87FDDF01FD0B33",
    X"FDDF01FD0B33FD1701D60B33",
    X"FF3503210F30FDDF03640F30",
    X"FDDF00000FADFF3503210F30",
    X"FF3503210F30FF2502FC0DFF",
    X"FF2502FC0DFFFDDF033C0DFF",
    X"FF2502FC0DFFFEA401CE0C87",
    X"FEA401CE0C87FDDF01F50C87",
    X"FEA401CE0C87FEA701D60B33",
    X"FEA701D60B33FDDF01FD0B33",
    X"004702690F30FF3503210F30",
    X"FDDF00000FAD004702690F30",
    X"004702690F30002B024C0DFF",
    X"002B024C0DFFFF2502FC0DFF",
    X"002B024C0DFFFF4301640C87",
    X"FF4301640C87FEA401CE0C87",
    X"FF4301640C87FF4901690B33",
    X"FF4901690B33FEA701D60B33",
    X"00FF01550F30004702690F30",
    X"FDDF00000FAD00FF01550F30",
    X"00FF01550F3000DA01450DFF",
    X"00DA01450DFF002B024C0DFF",
    X"00DA01450DFFFFAE00C50C87",
    X"FFAE00C50C87FF4301640C87",
    X"FFAE00C50C87FFB500C80B33",
    X"FFB500C80B33FF4901690B33",
    X"014200000F3000FF01550F30",
    X"011A00000DFF00DA01450DFF",
    X"FFD500000C87FFAE00C50C87",
    X"FFDD00000B33FFB500C80B33",
    X"FFB5FF380B33020FFE380A50",
    X"020FFE380A50026900000A50",
    X"026900000A50FFDD00000B33",
    X"020FFE380A500572FCC709B4",
    X"0572FCC709B40614000009B4",
    X"0614000009B4026900000A50",
    X"0572FCC709B4087CFB7C0919",
    X"087CFB7C0919096100000919",
    X"0961000009190614000009B4",
    X"087CFB7C091909CEFAEC0836",
    X"09CEFAEC08360ACF00000836",
    X"0ACF00000836096100000919",
    X"FF49FE970B330118FCC70A50",
    X"0118FCC70A50020FFE380A50",
    X"0118FCC70A5003B3FA2C09B4",
    X"03B3FA2C09B40572FCC709B4",
    X"03B3FA2C09B4060AF7D40919",
    X"060AF7D40919087CFB7C0919",
    X"060AF7D40919070EF6D00836",
    X"070EF6D0083609CEFAEC0836",
    X"FEA7FE2A0B33FFA7FBD00A50",
    X"FFA7FBD00A500118FCC70A50",
    X"FFA7FBD00A500117F86D09B4",
    X"0117F86D09B403B3FA2C09B4",
    X"0117F86D09B40263F5620919",
    X"0263F5620919060AF7D40919",
    X"0263F562091902F2F4100836",
    X"02F2F4100836070EF6D00836",
    X"FDDFFE030B33FDDFFB760A50",
    X"FDDFFB760A50FFA7FBD00A50",
    X"FDDFFB760A50FDDFF7CA09B4",
    X"FDDFF7CA09B40117F86D09B4",
    X"FDDFF7CA09B4FDDFF47E0919",
    X"FDDFF47E09190263F5620919",
    X"FDDFF47E0919FDDFF30F0836",
    X"FDDFF30F083602F2F4100836",
    X"FD17FE2A0B33FC17FBD00A50",
    X"FC17FBD00A50FDDFFB760A50",
    X"FC17FBD00A50FAA6F86D09B4",
    X"FAA6F86D09B4FDDFF7CA09B4",
    X"FAA6F86D09B4F95AF5620919",
    X"F95AF5620919FDDFF47E0919",
    X"F95AF5620919F8CBF4100836",
    X"F8CBF4100836FDDFF30F0836",
    X"FC75FE970B33FAA5FCC70A50",
    X"FAA5FCC70A50FC17FBD00A50",
    X"FAA5FCC70A50F80AFA2C09B4",
    X"F80AFA2C09B4FAA6F86D09B4",
    X"F80AFA2C09B4F5B3F7D40919",
    X"F5B3F7D40919F95AF5620919",
    X"F5B3F7D40919F4AFF6D00836",
    X"F4AFF6D00836F8CBF4100836",
    X"FC09FF380B33F9AEFE380A50",
    X"F9AEFE380A50FAA5FCC70A50",
    X"F9AEFE380A50F64BFCC709B4",
    X"F64BFCC709B4F80AFA2C09B4",
    X"F64BFCC709B4F341FB7C0919",
    X"F341FB7C0919F5B3F7D40919",
    X"F341FB7C0919F1EFFAEC0836",
    X"F1EFFAEC0836F4AFF6D00836",
    X"FBE100000B33F95400000A50",
    X"F95400000A50F9AEFE380A50",
    X"F95400000A50F5A8000009B4",
    X"F5A8000009B4F64BFCC709B4",
    X"F5A8000009B4F25C00000919",
    X"F25C00000919F341FB7C0919",
    X"F25C00000919F0EE00000836",
    X"F0EE00000836F1EFFAEC0836",
    X"FC0900C80B33F9AE01C80A50",
    X"F9AE01C80A50F95400000A50",
    X"F9AE01C80A50F64B033909B4",
    X"F64B033909B4F5A8000009B4",
    X"F64B033909B4F34104840919",
    X"F34104840919F25C00000919",
    X"F34104840919F1EF05140836",
    X"F1EF05140836F0EE00000836",
    X"FC7501690B33FAA503390A50",
    X"FAA503390A50F9AE01C80A50",
    X"FAA503390A50F80A05D409B4",
    X"F80A05D409B4F64B033909B4",
    X"F80A05D409B4F5B3082C0919",
    X"F5B3082C0919F34104840919",
    X"F5B3082C0919F4AF09300836",
    X"F4AF09300836F1EF05140836",
    X"FD1701D60B33FC1704300A50",
    X"FC1704300A50FAA503390A50",
    X"FC1704300A50FAA6079309B4",
    X"FAA6079309B4F80A05D409B4",
    X"FAA6079309B4F95A0A9E0919",
    X"F95A0A9E0919F5B3082C0919",
    X"F95A0A9E0919F8CB0BF00836",
    X"F8CB0BF00836F4AF09300836",
    X"FDDF01FD0B33FDDF048A0A50",
    X"FDDF048A0A50FC1704300A50",
    X"FDDF048A0A50FDDF083609B4",
    X"FDDF083609B4FAA6079309B4",
    X"FDDF083609B4FDDF0B820919",
    X"FDDF0B820919F95A0A9E0919",
    X"FDDF0B820919FDDF0CF10836",
    X"FDDF0CF10836F8CB0BF00836",
    X"FEA701D60B33FFA704300A50",
    X"FFA704300A50FDDF048A0A50",
    X"FFA704300A500117079309B4",
    X"0117079309B4FDDF083609B4",
    X"0117079309B402630A9E0919",
    X"02630A9E0919FDDF0B820919",
    X"02630A9E091902F20BF00836",
    X"02F20BF00836FDDF0CF10836",
    X"FF4901690B33011803390A50",
    X"011803390A50FFA704300A50",
    X"011803390A5003B305D409B4",
    X"03B305D409B40117079309B4",
    X"03B305D409B4060A082C0919",
    X"060A082C091902630A9E0919",
    X"060A082C0919070E09300836",
    X"070E0930083602F20BF00836",
    X"FFB500C80B33020F01C80A50",
    X"020F01C80A50011803390A50",
    X"020F01C80A500572033909B4",
    X"0572033909B403B305D409B4",
    X"0572033909B4087C04840919",
    X"087C04840919060A082C0919",
    X"087C0484091909CE05140836",
    X"09CE05140836070E09300836",
    X"026900000A50020F01C80A50",
    X"0614000009B40572033909B4",
    X"096100000919087C04840919",
    X"0ACF0000083609CE05140836"
  );
end package;